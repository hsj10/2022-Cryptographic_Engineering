`timescale 1ns/100ps 
module Key_Extension(input [64:1] key0,
				output reg [48:1] Key1, Key2, Key3, Key4, Key5, Key6, Key7, Key8, Key9, Key10, Key11, Key12, Key13, Key14, Key15, Key16);

  wire   [1:64] key;
  wire   [48:1] key1, key2, key3, key4, key5, key6, key7, key8, key9, key10, key11, key12, key13, key14, key15, key16;
  wire   [1:56] C0D0;
  wire   [1:56] C1D1;
  wire   [1:56] C2D2;
  wire   [1:56] C3D3;
  wire   [1:56] C4D4;
  wire   [1:56] C5D5;
  wire   [1:56] C6D6;
  wire   [1:56] C7D7;
  wire   [1:56] C8D8;
  wire   [1:56] C9D9;
  wire   [1:56] C10D10;
  wire   [1:56] C11D11;
  wire   [1:56] C12D12;
  wire   [1:56] C13D13;
  wire   [1:56] C14D14;
  wire   [1:56] C15D15;
  wire   [1:56] C16D16;


  assign key={key0[64],key0[63],key0[62],key0[61],key0[60],key0[59],key0[58],key0[57],key0[56],
  	key0[55],key0[54],key0[53],key0[52],key0[51],key0[50],key0[49],key0[48],key0[47],
  	key0[46],key0[45],key0[44],key0[43],key0[42],key0[41],key0[40],key0[39],key0[38],
  	key0[37],key0[36],key0[35],key0[34],key0[33],key0[32],key0[31],key0[30],key0[29],
  	key0[28],key0[27],key0[26],key0[25],key0[24],key0[23],key0[22],key0[21],key0[20],
  	key0[19],key0[18],key0[17],key0[16],key0[15],key0[14],key0[13],key0[12],key0[11],
  	key0[10],key0[9],key0[8],key0[7],key0[6],key0[5],key0[4],key0[3],key0[2],key0[1]};
  
  
  assign C0D0 = {
    key[57], key[49], key[41], key[33], key[25], key[17], key[09],
    key[01], key[58], key[50], key[42], key[34], key[26], key[18],
    key[10], key[02], key[59], key[51], key[43], key[35], key[27],
    key[19], key[11], key[03], key[60], key[52], key[44], key[36],
    key[63], key[55], key[47], key[39], key[31], key[23], key[15],
    key[07], key[62], key[54], key[46], key[38], key[30], key[22],
    key[14], key[06], key[61], key[53], key[45], key[37], key[29],
    key[21], key[13], key[05], key[28], key[20] ,key[12], key[04]
  };



  assign C1D1  = {C0D0[2:28],  C0D0[1],    C0D0[30:56],  C0D0[29]};
  assign C2D2  = {C1D1[2:28],  C1D1[1],    C1D1[30:56],  C1D1[29]};
  assign C3D3  = {C2D2[3:28],  C2D2[1:2],  C2D2[31:56],  C2D2[29:30]};
  assign C4D4  = {C3D3[3:28],  C3D3[1:2],  C3D3[31:56],  C3D3[29:30]};
  assign C5D5  = {C4D4[3:28],  C4D4[1:2],  C4D4[31:56],  C4D4[29:30]};
  assign C6D6  = {C5D5[3:28],  C5D5[1:2],  C5D5[31:56],  C5D5[29:30]};
  assign C7D7  = {C6D6[3:28],  C6D6[1:2],  C6D6[31:56],  C6D6[29:30]};
  assign C8D8  = {C7D7[3:28],  C7D7[1:2],  C7D7[31:56],  C7D7[29:30]};
  assign C9D9  = {C8D8[2:28],  C8D8[1],    C8D8[30:56],  C8D8[29]};
  assign C10D10= {C9D9[3:28],  C9D9[1:2],  C9D9[31:56],  C9D9[29:30]};
  assign C11D11= {C10D10[3:28],C10D10[1:2],C10D10[31:56],C10D10[29:30]};
  assign C12D12= {C11D11[3:28],C11D11[1:2],C11D11[31:56],C11D11[29:30]};
  assign C13D13= {C12D12[3:28],C12D12[1:2],C12D12[31:56],C12D12[29:30]};
  assign C14D14= {C13D13[3:28],C13D13[1:2],C13D13[31:56],C13D13[29:30]};
  assign C15D15= {C14D14[3:28],C14D14[1:2],C14D14[31:56],C14D14[29:30]};
  assign C16D16= {C15D15[2:28],C15D15[1],  C15D15[30:56],C15D15[29]};


  assign key1 = {
    C1D1[14],C1D1[17],C1D1[11],C1D1[24],C1D1[1], C1D1[5],
    C1D1[3] ,C1D1[28],C1D1[15],C1D1[6], C1D1[21],C1D1[10],
    C1D1[23],C1D1[19],C1D1[12],C1D1[4], C1D1[26],C1D1[8],
    C1D1[16],C1D1[7], C1D1[27],C1D1[20],C1D1[13],C1D1[2],
    C1D1[41],C1D1[52],C1D1[31],C1D1[37],C1D1[47],C1D1[55],
    C1D1[30],C1D1[40],C1D1[51],C1D1[45],C1D1[33],C1D1[48],
    C1D1[44],C1D1[49],C1D1[39],C1D1[56],C1D1[34],C1D1[53],
    C1D1[46],C1D1[42],C1D1[50],C1D1[36],C1D1[29],C1D1[32]
  };


  	assign key2 = {
C2D2[14],C2D2[17],C2D2[11],C2D2[24],C2D2[1], C2D2[5],
    C2D2[3] ,C2D2[28],C2D2[15],C2D2[6], C2D2[21],C2D2[10],
    C2D2[23],C2D2[19],C2D2[12],C2D2[4], C2D2[26],C2D2[8],
    C2D2[16],C2D2[7], C2D2[27],C2D2[20],C2D2[13],C2D2[2],
    C2D2[41],C2D2[52],C2D2[31],C2D2[37],C2D2[47],C2D2[55],
    C2D2[30],C2D2[40],C2D2[51],C2D2[45],C2D2[33],C2D2[48],
    C2D2[44],C2D2[49],C2D2[39],C2D2[56],C2D2[34],C2D2[53],
    C2D2[46],C2D2[42],C2D2[50],C2D2[36],C2D2[29],C2D2[32]
  };
  
	assign key3 = {
C3D3[14],C3D3[17],C3D3[11],C3D3[24],C3D3[1], C3D3[5],
    C3D3[3] ,C3D3[28],C3D3[15],C3D3[6], C3D3[21],C3D3[10],
    C3D3[23],C3D3[19],C3D3[12],C3D3[4], C3D3[26],C3D3[8],
    C3D3[16],C3D3[7], C3D3[27],C3D3[20],C3D3[13],C3D3[2],
    C3D3[41],C3D3[52],C3D3[31],C3D3[37],C3D3[47],C3D3[55],
    C3D3[30],C3D3[40],C3D3[51],C3D3[45],C3D3[33],C3D3[48],
    C3D3[44],C3D3[49],C3D3[39],C3D3[56],C3D3[34],C3D3[53],
    C3D3[46],C3D3[42],C3D3[50],C3D3[36],C3D3[29],C3D3[32]
  };

	assign key4 = {
C4D4[14],C4D4[17],C4D4[11],C4D4[24],C4D4[1], C4D4[5],
    C4D4[3] ,C4D4[28],C4D4[15],C4D4[6], C4D4[21],C4D4[10],
    C4D4[23],C4D4[19],C4D4[12],C4D4[4], C4D4[26],C4D4[8],
    C4D4[16],C4D4[7], C4D4[27],C4D4[20],C4D4[13],C4D4[2],
    C4D4[41],C4D4[52],C4D4[31],C4D4[37],C4D4[47],C4D4[55],
    C4D4[30],C4D4[40],C4D4[51],C4D4[45],C4D4[33],C4D4[48],
    C4D4[44],C4D4[49],C4D4[39],C4D4[56],C4D4[34],C4D4[53],
    C4D4[46],C4D4[42],C4D4[50],C4D4[36],C4D4[29],C4D4[32]
  };

	assign key5 = {
C5D5[14],C5D5[17],C5D5[11],C5D5[24],C5D5[1], C5D5[5],
    C5D5[3] ,C5D5[28],C5D5[15],C5D5[6], C5D5[21],C5D5[10],
    C5D5[23],C5D5[19],C5D5[12],C5D5[4], C5D5[26],C5D5[8],
    C5D5[16],C5D5[7], C5D5[27],C5D5[20],C5D5[13],C5D5[2],
    C5D5[41],C5D5[52],C5D5[31],C5D5[37],C5D5[47],C5D5[55],
    C5D5[30],C5D5[40],C5D5[51],C5D5[45],C5D5[33],C5D5[48],
    C5D5[44],C5D5[49],C5D5[39],C5D5[56],C5D5[34],C5D5[53],
    C5D5[46],C5D5[42],C5D5[50],C5D5[36],C5D5[29],C5D5[32]
  };
  	assign key6 = {
C6D6[14],C6D6[17],C6D6[11],C6D6[24],C6D6[1], C6D6[5],
    C6D6[3] ,C6D6[28],C6D6[15],C6D6[6], C6D6[21],C6D6[10],
    C6D6[23],C6D6[19],C6D6[12],C6D6[4], C6D6[26],C6D6[8],
    C6D6[16],C6D6[7], C6D6[27],C6D6[20],C6D6[13],C6D6[2],
    C6D6[41],C6D6[52],C6D6[31],C6D6[37],C6D6[47],C6D6[55],
    C6D6[30],C6D6[40],C6D6[51],C6D6[45],C6D6[33],C6D6[48],
    C6D6[44],C6D6[49],C6D6[39],C6D6[56],C6D6[34],C6D6[53],
    C6D6[46],C6D6[42],C6D6[50],C6D6[36],C6D6[29],C6D6[32]
  };

	assign key7 = {
C7D7[14],C7D7[17],C7D7[11],C7D7[24],C7D7[1], C7D7[5],
    C7D7[3] ,C7D7[28],C7D7[15],C7D7[6], C7D7[21],C7D7[10],
    C7D7[23],C7D7[19],C7D7[12],C7D7[4], C7D7[26],C7D7[8],
    C7D7[16],C7D7[7], C7D7[27],C7D7[20],C7D7[13],C7D7[2],
    C7D7[41],C7D7[52],C7D7[31],C7D7[37],C7D7[47],C7D7[55],
    C7D7[30],C7D7[40],C7D7[51],C7D7[45],C7D7[33],C7D7[48],
    C7D7[44],C7D7[49],C7D7[39],C7D7[56],C7D7[34],C7D7[53],
    C7D7[46],C7D7[42],C7D7[50],C7D7[36],C7D7[29],C7D7[32]
  };
	assign key8 = {
C8D8[14],C8D8[17],C8D8[11],C8D8[24],C8D8[1], C8D8[5],
    C8D8[3] ,C8D8[28],C8D8[15],C8D8[6], C8D8[21],C8D8[10],
    C8D8[23],C8D8[19],C8D8[12],C8D8[4], C8D8[26],C8D8[8],
    C8D8[16],C8D8[7], C8D8[27],C8D8[20],C8D8[13],C8D8[2],
    C8D8[41],C8D8[52],C8D8[31],C8D8[37],C8D8[47],C8D8[55],
    C8D8[30],C8D8[40],C8D8[51],C8D8[45],C8D8[33],C8D8[48],
    C8D8[44],C8D8[49],C8D8[39],C8D8[56],C8D8[34],C8D8[53],
    C8D8[46],C8D8[42],C8D8[50],C8D8[36],C8D8[29],C8D8[32]
  };
  
  	assign key9 = {
C9D9[14],C9D9[17],C9D9[11],C9D9[24],C9D9[1], C9D9[5],
    C9D9[3] ,C9D9[28],C9D9[15],C9D9[6], C9D9[21],C9D9[10],
    C9D9[23],C9D9[19],C9D9[12],C9D9[4], C9D9[26],C9D9[8],
    C9D9[16],C9D9[7], C9D9[27],C9D9[20],C9D9[13],C9D9[2],
    C9D9[41],C9D9[52],C9D9[31],C9D9[37],C9D9[47],C9D9[55],
    C9D9[30],C9D9[40],C9D9[51],C9D9[45],C9D9[33],C9D9[48],
    C9D9[44],C9D9[49],C9D9[39],C9D9[56],C9D9[34],C9D9[53],
    C9D9[46],C9D9[42],C9D9[50],C9D9[36],C9D9[29],C9D9[32]
  };
  
	assign key10 = {
C10D10[14],C10D10[17],C10D10[11],C10D10[24],C10D10[1], C10D10[5],
    C10D10[3] ,C10D10[28],C10D10[15],C10D10[6], C10D10[21],C10D10[10],
    C10D10[23],C10D10[19],C10D10[12],C10D10[4], C10D10[26],C10D10[8],
    C10D10[16],C10D10[7], C10D10[27],C10D10[20],C10D10[13],C10D10[2],
    C10D10[41],C10D10[52],C10D10[31],C10D10[37],C10D10[47],C10D10[55],
    C10D10[30],C10D10[40],C10D10[51],C10D10[45],C10D10[33],C10D10[48],
    C10D10[44],C10D10[49],C10D10[39],C10D10[56],C10D10[34],C10D10[53],
    C10D10[46],C10D10[42],C10D10[50],C10D10[36],C10D10[29],C10D10[32]
  };

	assign key11 = {
C11D11[14],C11D11[17],C11D11[11],C11D11[24],C11D11[1], C11D11[5],
    C11D11[3] ,C11D11[28],C11D11[15],C11D11[6], C11D11[21],C11D11[10],
    C11D11[23],C11D11[19],C11D11[12],C11D11[4], C11D11[26],C11D11[8],
    C11D11[16],C11D11[7], C11D11[27],C11D11[20],C11D11[13],C11D11[2],
    C11D11[41],C11D11[52],C11D11[31],C11D11[37],C11D11[47],C11D11[55],
    C11D11[30],C11D11[40],C11D11[51],C11D11[45],C11D11[33],C11D11[48],
    C11D11[44],C11D11[49],C11D11[39],C11D11[56],C11D11[34],C11D11[53],
    C11D11[46],C11D11[42],C11D11[50],C11D11[36],C11D11[29],C11D11[32]
  };

	assign key12 = {
C12D12[14],C12D12[17],C12D12[11],C12D12[24],C12D12[1], C12D12[5],
    C12D12[3] ,C12D12[28],C12D12[15],C12D12[6], C12D12[21],C12D12[10],
    C12D12[23],C12D12[19],C12D12[12],C12D12[4], C12D12[26],C12D12[8],
    C12D12[16],C12D12[7], C12D12[27],C12D12[20],C12D12[13],C12D12[2],
    C12D12[41],C12D12[52],C12D12[31],C12D12[37],C12D12[47],C12D12[55],
    C12D12[30],C12D12[40],C12D12[51],C12D12[45],C12D12[33],C12D12[48],
    C12D12[44],C12D12[49],C12D12[39],C12D12[56],C12D12[34],C12D12[53],
    C12D12[46],C12D12[42],C12D12[50],C12D12[36],C12D12[29],C12D12[32]
  };
  
  	assign key13 = {
C13D13[14],C13D13[17],C13D13[11],C13D13[24],C13D13[1], C13D13[5],
    C13D13[3] ,C13D13[28],C13D13[15],C13D13[6], C13D13[21],C13D13[10],
    C13D13[23],C13D13[19],C13D13[12],C13D13[4], C13D13[26],C13D13[8],
    C13D13[16],C13D13[7], C13D13[27],C13D13[20],C13D13[13],C13D13[2],
    C13D13[41],C13D13[52],C13D13[31],C13D13[37],C13D13[47],C13D13[55],
    C13D13[30],C13D13[40],C13D13[51],C13D13[45],C13D13[33],C13D13[48],
    C13D13[44],C13D13[49],C13D13[39],C13D13[56],C13D13[34],C13D13[53],
    C13D13[46],C13D13[42],C13D13[50],C13D13[36],C13D13[29],C13D13[32]
  };
  
	assign key14 = {
C14D14[14],C14D14[17],C14D14[11],C14D14[24],C14D14[1], C14D14[5],
    C14D14[3] ,C14D14[28],C14D14[15],C14D14[6], C14D14[21],C14D14[10],
    C14D14[23],C14D14[19],C14D14[12],C14D14[4], C14D14[26],C14D14[8],
    C14D14[16],C14D14[7], C14D14[27],C14D14[20],C14D14[13],C14D14[2],
    C14D14[41],C14D14[52],C14D14[31],C14D14[37],C14D14[47],C14D14[55],
    C14D14[30],C14D14[40],C14D14[51],C14D14[45],C14D14[33],C14D14[48],
    C14D14[44],C14D14[49],C14D14[39],C14D14[56],C14D14[34],C14D14[53],
    C14D14[46],C14D14[42],C14D14[50],C14D14[36],C14D14[29],C14D14[32]
  };
  
	assign key15 = {
C15D15[14],C15D15[17],C15D15[11],C15D15[24],C15D15[1], C15D15[5],
    C15D15[3] ,C15D15[28],C15D15[15],C15D15[6], C15D15[21],C15D15[10],
    C15D15[23],C15D15[19],C15D15[12],C15D15[4], C15D15[26],C15D15[8],
    C15D15[16],C15D15[7], C15D15[27],C15D15[20],C15D15[13],C15D15[2],
    C15D15[41],C15D15[52],C15D15[31],C15D15[37],C15D15[47],C15D15[55],
    C15D15[30],C15D15[40],C15D15[51],C15D15[45],C15D15[33],C15D15[48],
    C15D15[44],C15D15[49],C15D15[39],C15D15[56],C15D15[34],C15D15[53],
    C15D15[46],C15D15[42],C15D15[50],C15D15[36],C15D15[29],C15D15[32]
  };
  
	assign key16 = {
C16D16[14],C16D16[17],C16D16[11],C16D16[24],C16D16[1], C16D16[5],
    C16D16[3] ,C16D16[28],C16D16[15],C16D16[6], C16D16[21],C16D16[10],
    C16D16[23],C16D16[19],C16D16[12],C16D16[4], C16D16[26],C16D16[8],
    C16D16[16],C16D16[7], C16D16[27],C16D16[20],C16D16[13],C16D16[2],
    C16D16[41],C16D16[52],C16D16[31],C16D16[37],C16D16[47],C16D16[55],
    C16D16[30],C16D16[40],C16D16[51],C16D16[45],C16D16[33],C16D16[48],
    C16D16[44],C16D16[49],C16D16[39],C16D16[56],C16D16[34],C16D16[53],
    C16D16[46],C16D16[42],C16D16[50],C16D16[36],C16D16[29],C16D16[32]
  };
  
  always@(*)
  begin
  Key1<=key1;
  Key2<=key2;
  Key3<=key3;
  Key4<=key4;
  Key5<=key5;
  Key6<=key6;
  Key7<=key7;
  Key8<=key8;
  Key9<=key9;
  Key10<=key10;
  Key11<=key11;
  Key12<=key12;
  Key13<=key13;
  Key14<=key14;
  Key15<=key15;
  Key16<=key16;
end

//initial $monitor("Key1=%b,Key2=%b,Key3=%b,Key4=%b,Key5=%b,Key6=%b,Key7=%b,Key8=%b,Key9=%b,Key10=%b,Key11=%b,Key12=%b,Key13=%b,Key14=%b,Key15=%b,Key16=%b",Key1,Key2,Key3,Key4,Key5,Key6,Key7,Key8,Key9,Key10,Key11,Key12,Key13,Key14,Key15,Key16);


  
	endmodule
	
		
	
	